library verilog;
use verilog.vl_types.all;
entity \Chen_Kevin_SR-Latch\ is
    port(
        Chen_Kevin_Q    : out    vl_logic;
        Chen_Kevin_S    : in     vl_logic;
        Chen_Kevin_R    : in     vl_logic;
        Chen_Kevin_QNOT : out    vl_logic
    );
end \Chen_Kevin_SR-Latch\;
